`timescale 1ns / 1ps
module instRam(
        input pl_clk,
        input ps_clk,
        input [31:0] in_instruction,
        input [7:0] write_adr,
        input [7:0] read_adr,
        input w,
        input r,
        output reg [31:0] out_instruction, 
	    output [2:0] TMDSp, TMDSn,
	    output TMDSp_clock, TMDSn_clock
	   

    );
    reg [31:0] ram [255:0];
    wire [9:0] hdmi_x, hdmi_y;
    wire debiloba_r;
    wire [23:0] hdmi_c;
    wire [71:0] presents;
    
    always @(posedge ps_clk)
    begin
      
        
        if(w)
        begin
            ram[write_adr] <= in_instruction;
        end
        if(r)
        begin
            out_instruction <= ram[write_adr];
        end
    end
    
    HDMI_test(
	.clk(pl_clk),  // 125MHz
	//input valll,
	.vr(hdmi_c[7:0]),
	.vg(hdmi_c[15:8]),
	.vb(hdmi_c[23:16]),
	.TMDSp(TMDSp), .TMDSn(TMDSn),
	.TMDSp_clock(TMDSp_clock), .TMDSn_clock(TMDSn_clock),
	.xout(hdmi_x), .yout(hdmi_y),
	.r(debiloba_r)
    );
    
    assign hdmi_c = presents[0] ? ram[3][23:0] :
                presents[1] ? ram[7][23:0] :
                presents[2] ? ram[11][23:0] :
                presents[3] ? ram[15][23:0] :
                presents[4] ? ram[19][23:0] :
                presents[5] ? ram[23][23:0] :
                presents[6] ? ram[27][23:0] :
                presents[7] ? ram[31][23:0] :
                //circle
                presents[8] ? ram[33][23:0] :
                presents[9] ? ram[35][23:0] :
                presents[10] ? ram[37][23:0] :
                presents[11] ? ram[39][23:0] :
                presents[12] ? ram[41][23:0] :
                presents[13] ? ram[43][23:0] :
                presents[14] ? ram[45][23:0] :
                presents[15] ? ram[47][23:0] :
                presents[16] ? ram[49][23:0] :
                presents[17] ? ram[51][23:0] :
                presents[18] ? ram[53][23:0] :
                presents[19] ? ram[55][23:0] :
                presents[20] ? ram[57][23:0] :
                presents[21] ? ram[59][23:0] :
                presents[22] ? ram[61][23:0] :
                presents[23] ? ram[63][23:0] :
                presents[24] ? ram[65][23:0] :
                presents[25] ? ram[67][23:0] :
                presents[26] ? ram[69][23:0] :
                presents[27] ? ram[71][23:0] :
                presents[28] ? ram[73][23:0] :
                presents[29] ? ram[75][23:0] :
                presents[30] ? ram[77][23:0] :
                presents[31] ? ram[79][23:0] :
                presents[32] ? ram[81][23:0] :
                presents[33] ? ram[83][23:0] :
                presents[34] ? ram[85][23:0] :
                presents[35] ? ram[87][23:0] :
                presents[36] ? ram[89][23:0] :
                presents[37] ? ram[91][23:0] :
                presents[38] ? ram[93][23:0] :
                presents[39] ? ram[95][23:0] :
                //rect
                presents[40] ? ram[98][23:0] :
                presents[41] ? ram[101][23:0] :
                presents[42] ? ram[104][23:0] :
                presents[43] ? ram[107][23:0] :
                presents[44] ? ram[110][23:0] :
                presents[45] ? ram[113][23:0] :
                presents[46] ? ram[116][23:0] :
                presents[47] ? ram[119][23:0] :
                presents[48] ? ram[122][23:0] :
                presents[49] ? ram[125][23:0] :
                presents[50] ? ram[128][23:0] :
                presents[51] ? ram[131][23:0] :
                presents[52] ? ram[134][23:0] :
                presents[53] ? ram[137][23:0] :
                presents[54] ? ram[140][23:0] :
                presents[55] ? ram[143][23:0] :
                presents[56] ? ram[146][23:0] :
                presents[57] ? ram[149][23:0] :
                presents[58] ? ram[152][23:0] :
                presents[59] ? ram[155][23:0] :
                presents[60] ? ram[158][23:0] :
                presents[61] ? ram[161][23:0] :
                presents[62] ? ram[164][23:0] :
                presents[63] ? ram[167][23:0] :
                presents[64] ? ram[170][23:0] :
                presents[65] ? ram[173][23:0] :
                presents[66] ? ram[176][23:0] :
                presents[67] ? ram[179][23:0] :
                presents[68] ? ram[182][23:0] :
                presents[69] ? ram[185][23:0] :
                presents[70] ? ram[188][23:0] :
                presents[71] ? ram[191][23:0] :
                24'd0;
    
        is_in_triangle isintr0 (
                .vertex_1x(ram[0][9:0]), .vertex_1y(ram[0][19:10]),
                .vertex_2x(ram[1][9:0]), .vertex_2y(ram[1][19:10]),
                .vertex_3x(ram[2][9:0]), .vertex_3y(ram[2][19:10]),
                .x(hdmi_x), .y(hdmi_y),
                .present(presents[0]),
                .active(ram[3][24])
        );
        is_in_triangle isintr1 (
                .vertex_1x(ram[4][9:0]), .vertex_1y(ram[4][19:10]),
                .vertex_2x(ram[5][9:0]), .vertex_2y(ram[5][19:10]),
                .vertex_3x(ram[6][9:0]), .vertex_3y(ram[6][19:10]),
                .x(hdmi_x), .y(hdmi_y),
                .present(presents[1]),
                .active(ram[7][24])
        );
        is_in_triangle isintr2 (
                .vertex_1x(ram[8][9:0]), .vertex_1y(ram[8][19:10]),
                .vertex_2x(ram[9][9:0]), .vertex_2y(ram[9][19:10]),
                .vertex_3x(ram[10][9:0]), .vertex_3y(ram[10][19:10]),
                .x(hdmi_x), .y(hdmi_y),
                .present(presents[2]),
                .active(ram[11][24])
        );
        is_in_triangle isintr3 (
                .vertex_1x(ram[12][9:0]), .vertex_1y(ram[12][19:10]),
                .vertex_2x(ram[13][9:0]), .vertex_2y(ram[13][19:10]),
                .vertex_3x(ram[14][9:0]), .vertex_3y(ram[14][19:10]),
                .x(hdmi_x), .y(hdmi_y),
                .present(presents[3]),
                .active(ram[15][24])
        );
        is_in_triangle isintr4 (
                .vertex_1x(ram[16][9:0]), .vertex_1y(ram[16][19:10]),
                .vertex_2x(ram[17][9:0]), .vertex_2y(ram[17][19:10]),
                .vertex_3x(ram[18][9:0]), .vertex_3y(ram[18][19:10]),
                .x(hdmi_x), .y(hdmi_y),
                .present(presents[4]),
                .active(ram[19][24])
        );
        is_in_triangle isintr5 (
                .vertex_1x(ram[20][9:0]), .vertex_1y(ram[20][19:10]),
                .vertex_2x(ram[21][9:0]), .vertex_2y(ram[21][19:10]),
                .vertex_3x(ram[22][9:0]), .vertex_3y(ram[22][19:10]),
                .x(hdmi_x), .y(hdmi_y),
                .present(presents[5]),
                .active(ram[23][24])
        );
        is_in_triangle isintr6 (
                .vertex_1x(ram[24][9:0]), .vertex_1y(ram[24][19:10]),
                .vertex_2x(ram[25][9:0]), .vertex_2y(ram[25][19:10]),
                .vertex_3x(ram[26][9:0]), .vertex_3y(ram[26][19:10]),
                .x(hdmi_x), .y(hdmi_y),
                .present(presents[6]),
                .active(ram[27][24])
        );
        is_in_triangle isintr7 (
                .vertex_1x(ram[28][9:0]), .vertex_1y(ram[28][19:10]),
                .vertex_2x(ram[29][9:0]), .vertex_2y(ram[29][19:10]),
                .vertex_3x(ram[30][9:0]), .vertex_3y(ram[30][19:10]),
                .x(hdmi_x), .y(hdmi_y),
                .present(presents[7]),
                .active(ram[31][24])
        );
        in_circle c0(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[32][9:0]), .circle_y(ram[32][19:10]), .circle_rad(ram[32][29:20]),
                .active(ram[33][24]),
                .present(presents[8])
                );
        
        in_circle c1(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[34][9:0]), .circle_y(ram[34][19:10]), .circle_rad(ram[34][29:20]),
                .active(ram[35][24]),
                .present(presents[9])
                );
        
        in_circle c2(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[36][9:0]), .circle_y(ram[36][19:10]), .circle_rad(ram[36][29:20]),
                .active(ram[37][24]),
                .present(presents[10])
                );
        
        in_circle c3(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[38][9:0]), .circle_y(ram[38][19:10]), .circle_rad(ram[38][29:20]),
                .active(ram[39][24]),
                .present(presents[11])
                );
        
        in_circle c4(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[40][9:0]), .circle_y(ram[40][19:10]), .circle_rad(ram[40][29:20]),
                .active(ram[41][24]),
                .present(presents[12])
                );
        
        in_circle c5(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[42][9:0]), .circle_y(ram[42][19:10]), .circle_rad(ram[42][29:20]),
                .active(ram[43][24]),
                .present(presents[13])
                );
        
        in_circle c6(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[44][9:0]), .circle_y(ram[44][19:10]), .circle_rad(ram[44][29:20]),
                .active(ram[45][24]),
                .present(presents[14])
                );
        
        in_circle c7(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[46][9:0]), .circle_y(ram[46][19:10]), .circle_rad(ram[46][29:20]),
                .active(ram[47][24]),
                .present(presents[15])
                );
        
        in_circle c8(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[48][9:0]), .circle_y(ram[48][19:10]), .circle_rad(ram[48][29:20]),
                .active(ram[49][24]),
                .present(presents[16])
                );
        
        in_circle c9(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[50][9:0]), .circle_y(ram[50][19:10]), .circle_rad(ram[50][29:20]),
                .active(ram[51][24]),
                .present(presents[17])
                );
        
        in_circle c10(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[52][9:0]), .circle_y(ram[52][19:10]), .circle_rad(ram[52][29:20]),
                .active(ram[53][24]),
                .present(presents[18])
                );
        
        in_circle c11(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[54][9:0]), .circle_y(ram[54][19:10]), .circle_rad(ram[54][29:20]),
                .active(ram[55][24]),
                .present(presents[19])
                );
        
        in_circle c12(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[56][9:0]), .circle_y(ram[56][19:10]), .circle_rad(ram[56][29:20]),
                .active(ram[57][24]),
                .present(presents[20])
                );
        
        in_circle c13(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[58][9:0]), .circle_y(ram[58][19:10]), .circle_rad(ram[58][29:20]),
                .active(ram[59][24]),
                .present(presents[21])
                );
        
        in_circle c14(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[60][9:0]), .circle_y(ram[60][19:10]), .circle_rad(ram[60][29:20]),
                .active(ram[61][24]),
                .present(presents[22])
                );
        
        in_circle c15(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[62][9:0]), .circle_y(ram[62][19:10]), .circle_rad(ram[62][29:20]),
                .active(ram[63][24]),
                .present(presents[23])
                );
        
        in_circle c16(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[64][9:0]), .circle_y(ram[64][19:10]), .circle_rad(ram[64][29:20]),
                .active(ram[65][24]),
                .present(presents[24])
                );
        
        in_circle c17(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[66][9:0]), .circle_y(ram[66][19:10]), .circle_rad(ram[66][29:20]),
                .active(ram[67][24]),
                .present(presents[25])
                );
        
        in_circle c18(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[68][9:0]), .circle_y(ram[68][19:10]), .circle_rad(ram[68][29:20]),
                .active(ram[69][24]),
                .present(presents[26])
                );
        
        in_circle c19(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[70][9:0]), .circle_y(ram[70][19:10]), .circle_rad(ram[70][29:20]),
                .active(ram[71][24]),
                .present(presents[27])
                );
        
        in_circle c20(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[72][9:0]), .circle_y(ram[72][19:10]), .circle_rad(ram[72][29:20]),
                .active(ram[73][24]),
                .present(presents[28])
                );
        
        in_circle c21(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[74][9:0]), .circle_y(ram[74][19:10]), .circle_rad(ram[74][29:20]),
                .active(ram[75][24]),
                .present(presents[29])
                );
        
        in_circle c22(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[76][9:0]), .circle_y(ram[76][19:10]), .circle_rad(ram[76][29:20]),
                .active(ram[77][24]),
                .present(presents[30])
                );
        
        in_circle c23(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[78][9:0]), .circle_y(ram[78][19:10]), .circle_rad(ram[78][29:20]),
                .active(ram[79][24]),
                .present(presents[31])
                );
        
        in_circle c24(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[80][9:0]), .circle_y(ram[80][19:10]), .circle_rad(ram[80][29:20]),
                .active(ram[81][24]),
                .present(presents[32])
                );
        
        in_circle c25(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[82][9:0]), .circle_y(ram[82][19:10]), .circle_rad(ram[82][29:20]),
                .active(ram[83][24]),
                .present(presents[33])
                );
        
        in_circle c26(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[84][9:0]), .circle_y(ram[84][19:10]), .circle_rad(ram[84][29:20]),
                .active(ram[85][24]),
                .present(presents[34])
                );
        
        in_circle c27(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[86][9:0]), .circle_y(ram[86][19:10]), .circle_rad(ram[86][29:20]),
                .active(ram[87][24]),
                .present(presents[35])
                );
        
        in_circle c28(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[88][9:0]), .circle_y(ram[88][19:10]), .circle_rad(ram[88][29:20]),
                .active(ram[89][24]),
                .present(presents[36])
                );
        
        in_circle c29(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[90][9:0]), .circle_y(ram[90][19:10]), .circle_rad(ram[90][29:20]),
                .active(ram[91][24]),
                .present(presents[37])
                );
        
        in_circle c30(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[92][9:0]), .circle_y(ram[92][19:10]), .circle_rad(ram[92][29:20]),
                .active(ram[93][24]),
                .present(presents[38])
                );
        
        in_circle c31(
                .x(hdmi_x),.y(hdmi_y),
                .circle_x(ram[94][9:0]), .circle_y(ram[94][19:10]), .circle_rad(ram[94][29:20]),
                .active(ram[95][24]),
                .present(presents[39])
                );
        in_rect r0(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[96][9:0]), .rect_y(ram[96][19:10]), .rect_w(ram[97][9:0]), .rect_h(ram[97][19:10]),
                        .active(ram[98][24]),
                        .present(presents[40])
                        );
        in_rect r1(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[99][9:0]), .rect_y(ram[99][19:10]), .rect_w(ram[100][9:0]), .rect_h(ram[100][19:10]),
                        .active(ram[101][24]),
                        .present(presents[41])
                        );
        in_rect r2(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[102][9:0]), .rect_y(ram[102][19:10]), .rect_w(ram[103][9:0]), .rect_h(ram[103][19:10]),
                        .active(ram[104][24]),
                        .present(presents[42])
                        );
        in_rect r3(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[105][9:0]), .rect_y(ram[105][19:10]), .rect_w(ram[106][9:0]), .rect_h(ram[106][19:10]),
                        .active(ram[107][24]),
                        .present(presents[43])
                        );
        in_rect r4(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[108][9:0]), .rect_y(ram[108][19:10]), .rect_w(ram[109][9:0]), .rect_h(ram[109][19:10]),
                        .active(ram[110][24]),
                        .present(presents[44])
                        );
        in_rect r5(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[111][9:0]), .rect_y(ram[111][19:10]), .rect_w(ram[112][9:0]), .rect_h(ram[112][19:10]),
                        .active(ram[113][24]),
                        .present(presents[45])
                        );
        in_rect r6(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[114][9:0]), .rect_y(ram[114][19:10]), .rect_w(ram[115][9:0]), .rect_h(ram[115][19:10]),
                        .active(ram[116][24]),
                        .present(presents[46])
                        );
        in_rect r7(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[117][9:0]), .rect_y(ram[117][19:10]), .rect_w(ram[118][9:0]), .rect_h(ram[118][19:10]),
                        .active(ram[119][24]),
                        .present(presents[47])
                        );
        in_rect r8(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[120][9:0]), .rect_y(ram[120][19:10]), .rect_w(ram[121][9:0]), .rect_h(ram[121][19:10]),
                        .active(ram[122][24]),
                        .present(presents[48])
                        );
        in_rect r9(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[123][9:0]), .rect_y(ram[123][19:10]), .rect_w(ram[124][9:0]), .rect_h(ram[124][19:10]),
                        .active(ram[125][24]),
                        .present(presents[49])
                        );
        in_rect r10(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[126][9:0]), .rect_y(ram[126][19:10]), .rect_w(ram[127][9:0]), .rect_h(ram[127][19:10]),
                        .active(ram[128][24]),
                        .present(presents[50])
                        );
        in_rect r11(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[129][9:0]), .rect_y(ram[129][19:10]), .rect_w(ram[130][9:0]), .rect_h(ram[130][19:10]),
                        .active(ram[131][24]),
                        .present(presents[51])
                        );
        in_rect r12(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[132][9:0]), .rect_y(ram[132][19:10]), .rect_w(ram[133][9:0]), .rect_h(ram[133][19:10]),
                        .active(ram[134][24]),
                        .present(presents[52])
                        );
        in_rect r13(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[135][9:0]), .rect_y(ram[135][19:10]), .rect_w(ram[136][9:0]), .rect_h(ram[136][19:10]),
                        .active(ram[137][24]),
                        .present(presents[53])
                        );
        in_rect r14(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[138][9:0]), .rect_y(ram[138][19:10]), .rect_w(ram[139][9:0]), .rect_h(ram[139][19:10]),
                        .active(ram[140][24]),
                        .present(presents[54])
                        );
        in_rect r15(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[141][9:0]), .rect_y(ram[141][19:10]), .rect_w(ram[142][9:0]), .rect_h(ram[142][19:10]),
                        .active(ram[143][24]),
                        .present(presents[55])
                        );
        in_rect r16(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[144][9:0]), .rect_y(ram[144][19:10]), .rect_w(ram[145][9:0]), .rect_h(ram[145][19:10]),
                        .active(ram[146][24]),
                        .present(presents[56])
                        );
        in_rect r17(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[147][9:0]), .rect_y(ram[147][19:10]), .rect_w(ram[148][9:0]), .rect_h(ram[148][19:10]),
                        .active(ram[149][24]),
                        .present(presents[57])
                        );
        in_rect r18(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[150][9:0]), .rect_y(ram[150][19:10]), .rect_w(ram[151][9:0]), .rect_h(ram[151][19:10]),
                        .active(ram[152][24]),
                        .present(presents[58])
                        );
        in_rect r19(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[153][9:0]), .rect_y(ram[153][19:10]), .rect_w(ram[154][9:0]), .rect_h(ram[154][19:10]),
                        .active(ram[155][24]),
                        .present(presents[59])
                        );
        in_rect r20(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[156][9:0]), .rect_y(ram[156][19:10]), .rect_w(ram[157][9:0]), .rect_h(ram[157][19:10]),
                        .active(ram[158][24]),
                        .present(presents[60])
                        );
        in_rect r21(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[159][9:0]), .rect_y(ram[159][19:10]), .rect_w(ram[160][9:0]), .rect_h(ram[160][19:10]),
                        .active(ram[161][24]),
                        .present(presents[61])
                        );
        in_rect r22(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[162][9:0]), .rect_y(ram[162][19:10]), .rect_w(ram[163][9:0]), .rect_h(ram[163][19:10]),
                        .active(ram[164][24]),
                        .present(presents[62])
                        );
        in_rect r23(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[165][9:0]), .rect_y(ram[165][19:10]), .rect_w(ram[166][9:0]), .rect_h(ram[166][19:10]),
                        .active(ram[167][24]),
                        .present(presents[63])
                        );
        in_rect r24(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[168][9:0]), .rect_y(ram[168][19:10]), .rect_w(ram[169][9:0]), .rect_h(ram[169][19:10]),
                        .active(ram[170][24]),
                        .present(presents[64])
                        );
        in_rect r25(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[171][9:0]), .rect_y(ram[171][19:10]), .rect_w(ram[172][9:0]), .rect_h(ram[172][19:10]),
                        .active(ram[173][24]),
                        .present(presents[65])
                        );
        in_rect r26(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[174][9:0]), .rect_y(ram[174][19:10]), .rect_w(ram[175][9:0]), .rect_h(ram[175][19:10]),
                        .active(ram[176][24]),
                        .present(presents[66])
                        );
        in_rect r27(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[177][9:0]), .rect_y(ram[177][19:10]), .rect_w(ram[178][9:0]), .rect_h(ram[178][19:10]),
                        .active(ram[179][24]),
                        .present(presents[67])
                        );
        in_rect r28(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[180][9:0]), .rect_y(ram[180][19:10]), .rect_w(ram[181][9:0]), .rect_h(ram[181][19:10]),
                        .active(ram[182][24]),
                        .present(presents[68])
                        );
        in_rect r29(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[183][9:0]), .rect_y(ram[183][19:10]), .rect_w(ram[184][9:0]), .rect_h(ram[184][19:10]),
                        .active(ram[185][24]),
                        .present(presents[69])
                        );
        in_rect r30(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[186][9:0]), .rect_y(ram[186][19:10]), .rect_w(ram[187][9:0]), .rect_h(ram[187][19:10]),
                        .active(ram[188][24]),
                        .present(presents[70])
                        );
        in_rect r31(
                        .x(hdmi_x), .y(hdmi_y),
                        .rect_x(ram[189][9:0]), .rect_y(ram[189][19:10]), .rect_w(ram[190][9:0]), .rect_h(ram[190][19:10]),
                        .active(ram[191][24]),
                        .present(presents[71])
                        );
                
    
endmodule


